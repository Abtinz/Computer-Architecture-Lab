--------------------------------------------------------------------------------
-- Company: 
-- Engineer:
--
-- Create Date:   10:23:30 04/19/2022
-- Design Name:   
-- Module Name:   C:/Users/ABTIN/Documents/amirkabir un/term 4/Computer Architecture/Lab/HW6/RippleSubtractorAdder/TestBanch.vhd
-- Project Name:  RippleSubtractorAdder
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: FourBitRippleAdderSubtractor
-- 
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends
-- that these types always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--USE ieee.numeric_std.ALL;
 
ENTITY TestBanch IS
END TestBanch;
 
ARCHITECTURE behavior OF TestBanch IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT FourBitRippleAdderSubtractor
    PORT(
         A : IN  std_logic_vector(3 downto 0);
         B : IN  std_logic_vector(3 downto 0);
         Cin : IN  std_logic;
			Control_Signal : IN STD_LOGIC;
         Cout : OUT  std_logic;
         Sum : OUT  std_logic_vector(3 downto 0)
        );
    END COMPONENT;
    

   --Inputs
   signal A : std_logic_vector(3 downto 0) := (others => '0');
   signal B : std_logic_vector(3 downto 0) := (others => '0');
	signal Control_Signal : std_logic := '0';
   signal Cin : std_logic := '0';

 	--Outputs
   signal Cout : std_logic;
   signal Sum : std_logic_vector(3 downto 0);
   
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: FourBitRippleAdderSubtractor PORT MAP (
          A => A,
          B => B,
          Cin => Cin,
			 Control_Signal => Control_Signal ,
          Cout => Cout,
          Sum => Sum
        );


   stim_proc: process
   begin		
      -- hold reset state for 100 ns.
      wait for 100 ns;	

      A <= "1010";B<="1000"; Cin <= '0'; Control_Signal <= '0' ; wait for 100 ns;
		A <= "1110";B<="1001"; Cin <= '0'; Control_Signal <= '0' ; wait for 100 ns;
		A <= "1010";B<="1010"; Cin <= '0'; Control_Signal <= '0' ; wait for 100 ns;
		A <= "1001";B<="1110"; Cin <= '1'; Control_Signal <= '1' ; wait for 100 ns;
		A <= "1000";B<="1011"; Cin <= '1'; Control_Signal <= '1' ; wait for 100 ns;

      -- insert stimulus here 

      wait;
   end process;

END;
